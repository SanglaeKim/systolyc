// defines.sv --- 
// 
// Filename: defines.sv
// Description: 
// Author: Sanglae Kim
// Maintainer: 
// Created: Thu Dec 26 12:21:06 2024 (+0900)
// Version: 
// Package-Requires: ()
// Last-Updated: 
//           By: 
//     Update #: 0
// URL: 
// Doc URL: 
// Keywords: 
// Compatibility: 
// 
// 

// Code:
typedef struct{
   int pBase;
   int numBytes;
   string fileName;
}StSram;



// 
// defines.sv ends here
